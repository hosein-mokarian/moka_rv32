interface moka_rv32i_pipelined_if(input clk);
 logic rstn;
 logic en;
endinterface